library ieee;
use ieee.math_real.all;

package my_package is
	type dan_array is array (integer range 0 to 9 )
						of integer; -- lohlohloh
end my_package;